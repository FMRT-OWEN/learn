`include "./"
`include "./"

module ldst_select(
	)